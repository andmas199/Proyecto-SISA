LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE processor_components IS
    
END PACKAGE;