-- Listing 13.1
-- ROM with asynchonous read (inferring Block RAM)
-- character ROM
--   - 8-by-16 (8-by-2^4) font
--   - 256 (2^8) characters
--   - ROM size: 512-by-8 (2^11-by-8) bits
--               16K bits: 1 BRAM

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity vga_font_rom is
  port (
    clk  : in    std_logic;
    addr : in    std_logic_vector(11 downto 0);
    data : out   std_logic_vector(7 downto 0)
  );
end entity vga_font_rom;

architecture vga_font_rom_arch of vga_font_rom is

  constant addr_width : integer := 12;
  constant data_width : integer := 8;

  signal addr_reg : std_logic_vector(addr_width - 1 downto 0);

  type rom_type is array (0 to 2 ** addr_width - 1) of std_logic_vector(data_width - 1 downto 0);

  -- ROM definition
  constant rom : rom_type :=
  ( -- 2^11-by-8
    -- codigo x00
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x01
    "00000000", -- 0
    "00000000", -- 1
    "01111110", -- 2     ******
    "10000001", -- 3    *      *
    "10100101", -- 4    * *  * *
    "10000001", -- 5    *      *
    "10000001", -- 6    *      *
    "10111101", -- 7    * **** *
    "10011001", -- 8    *  **  *
    "10000001", -- 9    *      *
    "10000001", -- a    *      *
    "01111110", -- b     ******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x02
    "00000000", -- 0
    "00000000", -- 1
    "01111110", -- 2     ******
    "11111111", -- 3    ********
    "11011011", -- 4    ** ** **
    "11111111", -- 5    ********
    "11111111", -- 6    ********
    "11000011", -- 7    **    **
    "11100111", -- 8    ***  ***
    "11111111", -- 9    ********
    "11111111", -- a    ********
    "01111110", -- b     ******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x03
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "01101100", -- 4     ** **
    "11111110", -- 5    *******
    "11111110", -- 6    *******
    "11111110", -- 7    *******
    "11111110", -- 8    *******
    "01111100", -- 9     *****
    "00111000", -- a      ***
    "00010000", -- b       *
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x04
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00010000", -- 4       *
    "00111000", -- 5      ***
    "01111100", -- 6     *****
    "11111110", -- 7    *******
    "01111100", -- 8     *****
    "00111000", -- 9      ***
    "00010000", -- a       *
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x05
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00011000", -- 3       **
    "00111100", -- 4      ****
    "00111100", -- 5      ****
    "11100111", -- 6    ***  ***
    "11100111", -- 7    ***  ***
    "11100111", -- 8    ***  ***
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x06
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00011000", -- 3       **
    "00111100", -- 4      ****
    "01111110", -- 5     ******
    "11111111", -- 6    ********
    "11111111", -- 7    ********
    "01111110", -- 8     ******
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x07
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00011000", -- 6       **
    "00111100", -- 7      ****
    "00111100", -- 8      ****
    "00011000", -- 9       **
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x08
    "11111111", -- 0    ********
    "11111111", -- 1    ********
    "11111111", -- 2    ********
    "11111111", -- 3    ********
    "11111111", -- 4    ********
    "11111111", -- 5    ********
    "11100111", -- 6    ***  ***
    "11000011", -- 7    **    **
    "11000011", -- 8    **    **
    "11100111", -- 9    ***  ***
    "11111111", -- a    ********
    "11111111", -- b    ********
    "11111111", -- c    ********
    "11111111", -- d    ********
    "11111111", -- e    ********
    "11111111", -- f    ********
    -- codigo x09
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00111100", -- 5      ****
    "01100110", -- 6     **  **
    "01000010", -- 7     *    *
    "01000010", -- 8     *    *
    "01100110", -- 9     **  **
    "00111100", -- a      ****
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x0A
    "11111111", -- 0    ********
    "11111111", -- 1    ********
    "11111111", -- 2    ********
    "11111111", -- 3    ********
    "11111111", -- 4    ********
    "11000011", -- 5    **    **
    "10011001", -- 6    *  **  *
    "10111101", -- 7    * **** *
    "10111101", -- 8    * **** *
    "10011001", -- 9    *  **  *
    "11000011", -- a    **    **
    "11111111", -- b    ********
    "11111111", -- c    ********
    "11111111", -- d    ********
    "11111111", -- e    ********
    "11111111", -- f    ********
    -- codigo x0B
    "00000000", -- 0
    "00000000", -- 1
    "00011110", -- 2       ****
    "00001110", -- 3        ***
    "00011010", -- 4       ** *
    "00110010", -- 5      **  *
    "01111000", -- 6     ****
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01111000", -- b     ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x0C
    "00000000", -- 0
    "00000000", -- 1
    "00111100", -- 2      ****
    "01100110", -- 3     **  **
    "01100110", -- 4     **  **
    "01100110", -- 5     **  **
    "01100110", -- 6     **  **
    "00111100", -- 7      ****
    "00011000", -- 8       **
    "01111110", -- 9     ******
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x0D
    "00000000", -- 0
    "00000000", -- 1
    "00111111", -- 2      ******
    "00110011", -- 3      **  **
    "00111111", -- 4      ******
    "00110000", -- 5      **
    "00110000", -- 6      **
    "00110000", -- 7      **
    "00110000", -- 8      **
    "01110000", -- 9     ***
    "11110000", -- a    ****
    "11100000", -- b    ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x0E
    "00000000", -- 0
    "00000000", -- 1
    "01111111", -- 2     *******
    "01100011", -- 3     **   **
    "01111111", -- 4     *******
    "01100011", -- 5     **   **
    "01100011", -- 6     **   **
    "01100011", -- 7     **   **
    "01100011", -- 8     **   **
    "01100111", -- 9     **  ***
    "11100111", -- a    ***  ***
    "11100110", -- b    ***  **
    "11000000", -- c    **
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x0F
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00011000", -- 3       **
    "00011000", -- 4       **
    "11011011", -- 5    ** ** **
    "00111100", -- 6      ****
    "11100111", -- 7    ***  ***
    "00111100", -- 8      ****
    "11011011", -- 9    ** ** **
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x10
    "00000000", -- 0
    "10000000", -- 1    *
    "11000000", -- 2    **
    "11100000", -- 3    ***
    "11110000", -- 4    ****
    "11111000", -- 5    *****
    "11111110", -- 6    *******
    "11111000", -- 7    *****
    "11110000", -- 8    ****
    "11100000", -- 9    ***
    "11000000", -- a    **
    "10000000", -- b    *
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x11
    "00000000", -- 0
    "00000010", -- 1          *
    "00000110", -- 2         **
    "00001110", -- 3        ***
    "00011110", -- 4       ****
    "00111110", -- 5      *****
    "11111110", -- 6    *******
    "00111110", -- 7      *****
    "00011110", -- 8       ****
    "00001110", -- 9        ***
    "00000110", -- a         **
    "00000010", -- b          *
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x12
    "00000000", -- 0
    "00000000", -- 1
    "00011000", -- 2       **
    "00111100", -- 3      ****
    "01111110", -- 4     ******
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "01111110", -- 8     ******
    "00111100", -- 9      ****
    "00011000", -- a       **
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x13
    "00000000", -- 0
    "00000000", -- 1
    "01100110", -- 2     **  **
    "01100110", -- 3     **  **
    "01100110", -- 4     **  **
    "01100110", -- 5     **  **
    "01100110", -- 6     **  **
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "00000000", -- 9
    "01100110", -- a     **  **
    "01100110", -- b     **  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x14
    "00000000", -- 0
    "00000000", -- 1
    "01111111", -- 2     *******
    "11011011", -- 3    ** ** **
    "11011011", -- 4    ** ** **
    "11011011", -- 5    ** ** **
    "01111011", -- 6     **** **
    "00011011", -- 7       ** **
    "00011011", -- 8       ** **
    "00011011", -- 9       ** **
    "00011011", -- a       ** **
    "00011011", -- b       ** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x15
    "00000000", -- 0
    "01111100", -- 1     *****
    "11000110", -- 2    **   **
    "01100000", -- 3     **
    "00111000", -- 4      ***
    "01101100", -- 5     ** **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "01101100", -- 8     ** **
    "00111000", -- 9      ***
    "00001100", -- a        **
    "11000110", -- b    **   **
    "01111100", -- c     *****
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x16
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "11111110", -- 8    *******
    "11111110", -- 9    *******
    "11111110", -- a    *******
    "11111110", -- b    *******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x17
    "00000000", -- 0
    "00000000", -- 1
    "00011000", -- 2       **
    "00111100", -- 3      ****
    "01111110", -- 4     ******
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "01111110", -- 8     ******
    "00111100", -- 9      ****
    "00011000", -- a       **
    "01111110", -- b     ******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x18
    "00000000", -- 0
    "00000000", -- 1
    "00011000", -- 2       **
    "00111100", -- 3      ****
    "01111110", -- 4     ******
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x19
    "00000000", -- 0
    "00000000", -- 1
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "01111110", -- 9     ******
    "00111100", -- a      ****
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x1A
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00011000", -- 5       **
    "00001100", -- 6        **
    "11111110", -- 7    *******
    "00001100", -- 8        **
    "00011000", -- 9       **
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x1B
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00110000", -- 5      **
    "01100000", -- 6     **
    "11111110", -- 7    *******
    "01100000", -- 8     **
    "00110000", -- 9      **
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x1C
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "11000000", -- 6    **
    "11000000", -- 7    **
    "11000000", -- 8    **
    "11111110", -- 9    *******
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x1D
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00100100", -- 5      *  *
    "01100110", -- 6     **  **
    "11111111", -- 7    ********
    "01100110", -- 8     **  **
    "00100100", -- 9      *  *
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x1E
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00010000", -- 4       *
    "00111000", -- 5      ***
    "00111000", -- 6      ***
    "01111100", -- 7     *****
    "01111100", -- 8     *****
    "11111110", -- 9    *******
    "11111110", -- a    *******
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x1F
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "11111110", -- 4    *******
    "11111110", -- 5    *******
    "01111100", -- 6     *****
    "01111100", -- 7     *****
    "00111000", -- 8      ***
    "00111000", -- 9      ***
    "00010000", -- a       *
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x20
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x21
    "00000000", -- 0
    "00000000", -- 1
    "00011000", -- 2       **
    "00111100", -- 3      ****
    "00111100", -- 4      ****
    "00111100", -- 5      ****
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00000000", -- 9
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x22
    "00000000", -- 0
    "01100110", -- 1     **  **
    "01100110", -- 2     **  **
    "01100110", -- 3     **  **
    "00100100", -- 4      *  *
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x23
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "01101100", -- 3     ** **
    "01101100", -- 4     ** **
    "11111110", -- 5    *******
    "01101100", -- 6     ** **
    "01101100", -- 7     ** **
    "01101100", -- 8     ** **
    "11111110", -- 9    *******
    "01101100", -- a     ** **
    "01101100", -- b     ** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x24
    "00011000", -- 0       **
    "00011000", -- 1       **
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "11000010", -- 4    **    *
    "11000000", -- 5    **
    "01111100", -- 6     *****
    "00000110", -- 7         **
    "00000110", -- 8         **
    "10000110", -- 9    *    **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00011000", -- c       **
    "00011000", -- d       **
    "00000000", -- e
    "00000000", -- f
    -- codigo x25
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "11000010", -- 4    **    *
    "11000110", -- 5    **   **
    "00001100", -- 6        **
    "00011000", -- 7       **
    "00110000", -- 8      **
    "01100000", -- 9     **
    "11000110", -- a    **   **
    "10000110", -- b    *    **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x26
    "00000000", -- 0
    "00000000", -- 1
    "00111000", -- 2      ***
    "01101100", -- 3     ** **
    "01101100", -- 4     ** **
    "00111000", -- 5      ***
    "01110110", -- 6     *** **
    "11011100", -- 7    ** ***
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x27
    "00000000", -- 0
    "00110000", -- 1      **
    "00110000", -- 2      **
    "00110000", -- 3      **
    "01100000", -- 4     **
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x28
    "00000000", -- 0
    "00000000", -- 1
    "00001100", -- 2        **
    "00011000", -- 3       **
    "00110000", -- 4      **
    "00110000", -- 5      **
    "00110000", -- 6      **
    "00110000", -- 7      **
    "00110000", -- 8      **
    "00110000", -- 9      **
    "00011000", -- a       **
    "00001100", -- b        **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x29
    "00000000", -- 0
    "00000000", -- 1
    "00110000", -- 2      **
    "00011000", -- 3       **
    "00001100", -- 4        **
    "00001100", -- 5        **
    "00001100", -- 6        **
    "00001100", -- 7        **
    "00001100", -- 8        **
    "00001100", -- 9        **
    "00011000", -- a       **
    "00110000", -- b      **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x2A
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01100110", -- 5     **  **
    "00111100", -- 6      ****
    "11111111", -- 7    ********
    "00111100", -- 8      ****
    "01100110", -- 9     **  **
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x2B
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00011000", -- 5       **
    "00011000", -- 6       **
    "01111110", -- 7     ******
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x2C
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00110000", -- c      **
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x2D
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "11111110", -- 7    *******
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x2E
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x2Ff
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000010", -- 4          *
    "00000110", -- 5         **
    "00001100", -- 6        **
    "00011000", -- 7       **
    "00110000", -- 8      **
    "01100000", -- 9     **
    "11000000", -- a    **
    "10000000", -- b    *
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x30
    "00000000", -- 0
    "00000000", -- 1
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "11001110", -- 5    **  ***
    "11011110", -- 6    ** ****
    "11110110", -- 7    **** **
    "11100110", -- 8    ***  **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x31
    "00000000", -- 0
    "00000000", -- 1
    "00011000", -- 2       **
    "00111000", -- 3      ***
    "01111000", -- 4     ****
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "01111110", -- b     ******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x32
    "00000000", -- 0
    "00000000", -- 1
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "00000110", -- 4         **
    "00001100", -- 5        **
    "00011000", -- 6       **
    "00110000", -- 7      **
    "01100000", -- 8     **
    "11000000", -- 9    **
    "11000110", -- a    **   **
    "11111110", -- b    *******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x33
    "00000000", -- 0
    "00000000", -- 1
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "00000110", -- 4         **
    "00000110", -- 5         **
    "00111100", -- 6      ****
    "00000110", -- 7         **
    "00000110", -- 8         **
    "00000110", -- 9         **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x34
    "00000000", -- 0
    "00000000", -- 1
    "00001100", -- 2        **
    "00011100", -- 3       ***
    "00111100", -- 4      ****
    "01101100", -- 5     ** **
    "11001100", -- 6    **  **
    "11111110", -- 7    *******
    "00001100", -- 8        **
    "00001100", -- 9        **
    "00001100", -- a        **
    "00011110", -- b       ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x35
    "00000000", -- 0
    "00000000", -- 1
    "11111110", -- 2    *******
    "11000000", -- 3    **
    "11000000", -- 4    **
    "11000000", -- 5    **
    "11111100", -- 6    ******
    "00000110", -- 7         **
    "00000110", -- 8         **
    "00000110", -- 9         **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x36
    "00000000", -- 0
    "00000000", -- 1
    "00111000", -- 2      ***
    "01100000", -- 3     **
    "11000000", -- 4    **
    "11000000", -- 5    **
    "11111100", -- 6    ******
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x37
    "00000000", -- 0
    "00000000", -- 1
    "11111110", -- 2    *******
    "11000110", -- 3    **   **
    "00000110", -- 4         **
    "00000110", -- 5         **
    "00001100", -- 6        **
    "00011000", -- 7       **
    "00110000", -- 8      **
    "00110000", -- 9      **
    "00110000", -- a      **
    "00110000", -- b      **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x38
    "00000000", -- 0
    "00000000", -- 1
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "01111100", -- 6     *****
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x39
    "00000000", -- 0
    "00000000", -- 1
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "01111110", -- 6     ******
    "00000110", -- 7         **
    "00000110", -- 8         **
    "00000110", -- 9         **
    "00001100", -- a        **
    "01111000", -- b     ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x3A
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00011000", -- 9       **
    "00011000", -- a       **
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x3B
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00011000", -- 9       **
    "00011000", -- a       **
    "00110000", -- b      **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x3C
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000110", -- 3         **
    "00001100", -- 4        **
    "00011000", -- 5       **
    "00110000", -- 6      **
    "01100000", -- 7     **
    "00110000", -- 8      **
    "00011000", -- 9       **
    "00001100", -- a        **
    "00000110", -- b         **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x3D
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01111110", -- 5     ******
    "00000000", -- 6
    "00000000", -- 7
    "01111110", -- 8     ******
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x3E
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "01100000", -- 3     **
    "00110000", -- 4      **
    "00011000", -- 5       **
    "00001100", -- 6        **
    "00000110", -- 7         **
    "00001100", -- 8        **
    "00011000", -- 9       **
    "00110000", -- a      **
    "01100000", -- b     **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x3F
    "00000000", -- 0
    "00000000", -- 1
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "00001100", -- 5        **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00000000", -- 9
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x40
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "01111100", -- 3     *****
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "11011110", -- 6    ** ****
    "11011110", -- 7    ** ****
    "11011110", -- 8    ** ****
    "11011100", -- 9    ** ***
    "11000000", -- a    **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x41
    "00000000", -- 0
    "00000000", -- 1
    "00010000", -- 2       *
    "00111000", -- 3      ***
    "01101100", -- 4     ** **
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11111110", -- 7    *******
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "11000110", -- b    **   **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x42
    "00000000", -- 0
    "00000000", -- 1
    "11111100", -- 2    ******
    "01100110", -- 3     **  **
    "01100110", -- 4     **  **
    "01100110", -- 5     **  **
    "01111100", -- 6     *****
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "11111100", -- b    ******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x43
    "00000000", -- 0
    "00000000", -- 1
    "00111100", -- 2      ****
    "01100110", -- 3     **  **
    "11000010", -- 4    **    *
    "11000000", -- 5    **
    "11000000", -- 6    **
    "11000000", -- 7    **
    "11000000", -- 8    **
    "11000010", -- 9    **    *
    "01100110", -- a     **  **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x44
    "00000000", -- 0
    "00000000", -- 1
    "11111000", -- 2    *****
    "01101100", -- 3     ** **
    "01100110", -- 4     **  **
    "01100110", -- 5     **  **
    "01100110", -- 6     **  **
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01101100", -- a     ** **
    "11111000", -- b    *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x45
    "00000000", -- 0
    "00000000", -- 1
    "11111110", -- 2    *******
    "01100110", -- 3     **  **
    "01100010", -- 4     **   *
    "01101000", -- 5     ** *
    "01111000", -- 6     ****
    "01101000", -- 7     ** *
    "01100000", -- 8     **
    "01100010", -- 9     **   *
    "01100110", -- a     **  **
    "11111110", -- b    *******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x46
    "00000000", -- 0
    "00000000", -- 1
    "11111110", -- 2    *******
    "01100110", -- 3     **  **
    "01100010", -- 4     **   *
    "01101000", -- 5     ** *
    "01111000", -- 6     ****
    "01101000", -- 7     ** *
    "01100000", -- 8     **
    "01100000", -- 9     **
    "01100000", -- a     **
    "11110000", -- b    ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x47
    "00000000", -- 0
    "00000000", -- 1
    "00111100", -- 2      ****
    "01100110", -- 3     **  **
    "11000010", -- 4    **    *
    "11000000", -- 5    **
    "11000000", -- 6    **
    "11011110", -- 7    ** ****
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "01100110", -- a     **  **
    "00111010", -- b      *** *
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x48
    "00000000", -- 0
    "00000000", -- 1
    "11000110", -- 2    **   **
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "11111110", -- 6    *******
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "11000110", -- b    **   **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x49
    "00000000", -- 0
    "00000000", -- 1
    "00111100", -- 2      ****
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x4A
    "00000000", -- 0
    "00000000", -- 1
    "00011110", -- 2       ****
    "00001100", -- 3        **
    "00001100", -- 4        **
    "00001100", -- 5        **
    "00001100", -- 6        **
    "00001100", -- 7        **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01111000", -- b     ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x4B
    "00000000", -- 0
    "00000000", -- 1
    "11100110", -- 2    ***  **
    "01100110", -- 3     **  **
    "01100110", -- 4     **  **
    "01101100", -- 5     ** **
    "01111000", -- 6     ****
    "01111000", -- 7     ****
    "01101100", -- 8     ** **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "11100110", -- b    ***  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x4C
    "00000000", -- 0
    "00000000", -- 1
    "11110000", -- 2    ****
    "01100000", -- 3     **
    "01100000", -- 4     **
    "01100000", -- 5     **
    "01100000", -- 6     **
    "01100000", -- 7     **
    "01100000", -- 8     **
    "01100010", -- 9     **   *
    "01100110", -- a     **  **
    "11111110", -- b    *******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x4D
    "00000000", -- 0
    "00000000", -- 1
    "11000011", -- 2    **    **
    "11100111", -- 3    ***  ***
    "11111111", -- 4    ********
    "11111111", -- 5    ********
    "11011011", -- 6    ** ** **
    "11000011", -- 7    **    **
    "11000011", -- 8    **    **
    "11000011", -- 9    **    **
    "11000011", -- a    **    **
    "11000011", -- b    **    **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x4E
    "00000000", -- 0
    "00000000", -- 1
    "11000110", -- 2    **   **
    "11100110", -- 3    ***  **
    "11110110", -- 4    **** **
    "11111110", -- 5    *******
    "11011110", -- 6    ** ****
    "11001110", -- 7    **  ***
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "11000110", -- b    **   **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x4F
    "00000000", -- 0
    "00000000", -- 1
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x50
    "00000000", -- 0
    "00000000", -- 1
    "11111100", -- 2    ******
    "01100110", -- 3     **  **
    "01100110", -- 4     **  **
    "01100110", -- 5     **  **
    "01111100", -- 6     *****
    "01100000", -- 7     **
    "01100000", -- 8     **
    "01100000", -- 9     **
    "01100000", -- a     **
    "11110000", -- b    ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x51
    "00000000", -- 0
    "00000000", -- 1
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11010110", -- 9    ** * **
    "11011110", -- a    ** ****
    "01111100", -- b     *****
    "00001100", -- c        **
    "00001110", -- d        ***
    "00000000", -- e
    "00000000", -- f
    -- codigo x52
    "00000000", -- 0
    "00000000", -- 1
    "11111100", -- 2    ******
    "01100110", -- 3     **  **
    "01100110", -- 4     **  **
    "01100110", -- 5     **  **
    "01111100", -- 6     *****
    "01101100", -- 7     ** **
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "11100110", -- b    ***  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x53
    "00000000", -- 0
    "00000000", -- 1
    "01111100", -- 2     *****
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "01100000", -- 5     **
    "00111000", -- 6      ***
    "00001100", -- 7        **
    "00000110", -- 8         **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x54
    "00000000", -- 0
    "00000000", -- 1
    "11111111", -- 2    ********
    "11011011", -- 3    ** ** **
    "10011001", -- 4    *  **  *
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x55
    "00000000", -- 0
    "00000000", -- 1
    "11000110", -- 2    **   **
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x56
    "00000000", -- 0
    "00000000", -- 1
    "11000011", -- 2    **    **
    "11000011", -- 3    **    **
    "11000011", -- 4    **    **
    "11000011", -- 5    **    **
    "11000011", -- 6    **    **
    "11000011", -- 7    **    **
    "11000011", -- 8    **    **
    "01100110", -- 9     **  **
    "00111100", -- a      ****
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x57
    "00000000", -- 0
    "00000000", -- 1
    "11000011", -- 2    **    **
    "11000011", -- 3    **    **
    "11000011", -- 4    **    **
    "11000011", -- 5    **    **
    "11000011", -- 6    **    **
    "11011011", -- 7    ** ** **
    "11011011", -- 8    ** ** **
    "11111111", -- 9    ********
    "01100110", -- a     **  **
    "01100110", -- b     **  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x58
    "00000000", -- 0
    "00000000", -- 1
    "11000011", -- 2    **    **
    "11000011", -- 3    **    **
    "01100110", -- 4     **  **
    "00111100", -- 5      ****
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00111100", -- 8      ****
    "01100110", -- 9     **  **
    "11000011", -- a    **    **
    "11000011", -- b    **    **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x59
    "00000000", -- 0
    "00000000", -- 1
    "11000011", -- 2    **    **
    "11000011", -- 3    **    **
    "11000011", -- 4    **    **
    "01100110", -- 5     **  **
    "00111100", -- 6      ****
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x5A
    "00000000", -- 0
    "00000000", -- 1
    "11111111", -- 2    ********
    "11000011", -- 3    **    **
    "10000110", -- 4    *    **
    "00001100", -- 5        **
    "00011000", -- 6       **
    "00110000", -- 7      **
    "01100000", -- 8     **
    "11000001", -- 9    **     *
    "11000011", -- a    **    **
    "11111111", -- b    ********
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x5B
    "00000000", -- 0
    "00000000", -- 1
    "00111100", -- 2      ****
    "00110000", -- 3      **
    "00110000", -- 4      **
    "00110000", -- 5      **
    "00110000", -- 6      **
    "00110000", -- 7      **
    "00110000", -- 8      **
    "00110000", -- 9      **
    "00110000", -- a      **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x5C
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "10000000", -- 3    *
    "11000000", -- 4    **
    "11100000", -- 5    ***
    "01110000", -- 6     ***
    "00111000", -- 7      ***
    "00011100", -- 8       ***
    "00001110", -- 9        ***
    "00000110", -- a         **
    "00000010", -- b          *
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x5D
    "00000000", -- 0
    "00000000", -- 1
    "00111100", -- 2      ****
    "00001100", -- 3        **
    "00001100", -- 4        **
    "00001100", -- 5        **
    "00001100", -- 6        **
    "00001100", -- 7        **
    "00001100", -- 8        **
    "00001100", -- 9        **
    "00001100", -- a        **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x5E
    "00010000", -- 0       *
    "00111000", -- 1      ***
    "01101100", -- 2     ** **
    "11000110", -- 3    **   **
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x5F
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "11111111", -- d    ********
    "00000000", -- e
    "00000000", -- f
    -- codigo x60
    "00110000", -- 0      **
    "00110000", -- 1      **
    "00011000", -- 2       **
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x61
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01111000", -- 5     ****
    "00001100", -- 6        **
    "01111100", -- 7     *****
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x62
    "00000000", -- 0
    "00000000", -- 1
    "11100000", -- 2    ***
    "01100000", -- 3     **
    "01100000", -- 4     **
    "01111000", -- 5     ****
    "01101100", -- 6     ** **
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x63
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11000000", -- 7    **
    "11000000", -- 8    **
    "11000000", -- 9    **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x64
    "00000000", -- 0
    "00000000", -- 1
    "00011100", -- 2       ***
    "00001100", -- 3        **
    "00001100", -- 4        **
    "00111100", -- 5      ****
    "01101100", -- 6     ** **
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x65
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11111110", -- 7    *******
    "11000000", -- 8    **
    "11000000", -- 9    **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x66
    "00000000", -- 0
    "00000000", -- 1
    "00111000", -- 2      ***
    "01101100", -- 3     ** **
    "01100100", -- 4     **  *
    "01100000", -- 5     **
    "11110000", -- 6    ****
    "01100000", -- 7     **
    "01100000", -- 8     **
    "01100000", -- 9     **
    "01100000", -- a     **
    "11110000", -- b    ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x67
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01110110", -- 5     *** **
    "11001100", -- 6    **  **
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01111100", -- b     *****
    "00001100", -- c        **
    "11001100", -- d    **  **
    "01111000", -- e     ****
    "00000000", -- f
    -- codigo x68
    "00000000", -- 0
    "00000000", -- 1
    "11100000", -- 2    ***
    "01100000", -- 3     **
    "01100000", -- 4     **
    "01101100", -- 5     ** **
    "01110110", -- 6     *** **
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "11100110", -- b    ***  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x69
    "00000000", -- 0
    "00000000", -- 1
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00000000", -- 4
    "00111000", -- 5      ***
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x6A
    "00000000", -- 0
    "00000000", -- 1
    "00000110", -- 2         **
    "00000110", -- 3         **
    "00000000", -- 4
    "00001110", -- 5        ***
    "00000110", -- 6         **
    "00000110", -- 7         **
    "00000110", -- 8         **
    "00000110", -- 9         **
    "00000110", -- a         **
    "00000110", -- b         **
    "01100110", -- c     **  **
    "01100110", -- d     **  **
    "00111100", -- e      ****
    "00000000", -- f
    -- codigo x6B
    "00000000", -- 0
    "00000000", -- 1
    "11100000", -- 2    ***
    "01100000", -- 3     **
    "01100000", -- 4     **
    "01100110", -- 5     **  **
    "01101100", -- 6     ** **
    "01111000", -- 7     ****
    "01111000", -- 8     ****
    "01101100", -- 9     ** **
    "01100110", -- a     **  **
    "11100110", -- b    ***  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x6C
    "00000000", -- 0
    "00000000", -- 1
    "00111000", -- 2      ***
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x6D
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11100110", -- 5    ***  **
    "11111111", -- 6    ********
    "11011011", -- 7    ** ** **
    "11011011", -- 8    ** ** **
    "11011011", -- 9    ** ** **
    "11011011", -- a    ** ** **
    "11011011", -- b    ** ** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x6E
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11011100", -- 5    ** ***
    "01100110", -- 6     **  **
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "01100110", -- b     **  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x6F
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x70
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11011100", -- 5    ** ***
    "01100110", -- 6     **  **
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "01111100", -- b     *****
    "01100000", -- c     **
    "01100000", -- d     **
    "11110000", -- e    ****
    "00000000", -- f
    -- codigo x71
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01110110", -- 5     *** **
    "11001100", -- 6    **  **
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01111100", -- b     *****
    "00001100", -- c        **
    "00001100", -- d        **
    "00011110", -- e       ****
    "00000000", -- f
    -- codigo x72
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11011100", -- 5    ** ***
    "01110110", -- 6     *** **
    "01100110", -- 7     **  **
    "01100000", -- 8     **
    "01100000", -- 9     **
    "01100000", -- a     **
    "11110000", -- b    ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x73
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "01100000", -- 7     **
    "00111000", -- 8      ***
    "00001100", -- 9        **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x74
    "00000000", -- 0
    "00000000", -- 1
    "00010000", -- 2       *
    "00110000", -- 3      **
    "00110000", -- 4      **
    "11111100", -- 5    ******
    "00110000", -- 6      **
    "00110000", -- 7      **
    "00110000", -- 8      **
    "00110000", -- 9      **
    "00110110", -- a      ** **
    "00011100", -- b       ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x75
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11001100", -- 5    **  **
    "11001100", -- 6    **  **
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x76
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11000011", -- 5    **    **
    "11000011", -- 6    **    **
    "11000011", -- 7    **    **
    "11000011", -- 8    **    **
    "01100110", -- 9     **  **
    "00111100", -- a      ****
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x77
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11000011", -- 5    **    **
    "11000011", -- 6    **    **
    "11000011", -- 7    **    **
    "11011011", -- 8    ** ** **
    "11011011", -- 9    ** ** **
    "11111111", -- a    ********
    "01100110", -- b     **  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x78
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11000011", -- 5    **    **
    "01100110", -- 6     **  **
    "00111100", -- 7      ****
    "00011000", -- 8       **
    "00111100", -- 9      ****
    "01100110", -- a     **  **
    "11000011", -- b    **    **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x79
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111110", -- b     ******
    "00000110", -- c         **
    "00001100", -- d        **
    "11111000", -- e    *****
    "00000000", -- f
    -- codigo x7A
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11111110", -- 5    *******
    "11001100", -- 6    **  **
    "00011000", -- 7       **
    "00110000", -- 8      **
    "01100000", -- 9     **
    "11000110", -- a    **   **
    "11111110", -- b    *******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x7B
    "00000000", -- 0
    "00000000", -- 1
    "00001110", -- 2        ***
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "01110000", -- 6     ***
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00001110", -- b        ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x7C
    "00000000", -- 0
    "00000000", -- 1
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00000000", -- 6
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x7D
    "00000000", -- 0
    "00000000", -- 1
    "01110000", -- 2     ***
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00001110", -- 6        ***
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "01110000", -- b     ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x7E
    "00000000", -- 0
    "00000000", -- 1
    "01110110", -- 2     *** **
    "11011100", -- 3    ** ***
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x7Ff
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00010000", -- 4       *
    "00111000", -- 5      ***
    "01101100", -- 6     ** **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11111110", -- a    *******
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x80
    "00000000", -- 0
    "00000000", -- 1
    "00111100", -- 2      ****
    "01100110", -- 3     **  **
    "11000010", -- 4    **    *
    "11000000", -- 5    **
    "11000000", -- 6    **
    "11000000", -- 7    **
    "11000010", -- 8    **    *
    "01100110", -- 9     **  **
    "00111100", -- a      ****
    "00001100", -- b        **
    "00000110", -- c         **
    "01111100", -- d     *****
    "00000000", -- e
    "00000000", -- f
    -- codigo x81
    "00000000", -- 0
    "00000000", -- 1
    "11001100", -- 2    **  **
    "00000000", -- 3
    "00000000", -- 4
    "11001100", -- 5    **  **
    "11001100", -- 6    **  **
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x82
    "00000000", -- 0
    "00001100", -- 1        **
    "00011000", -- 2       **
    "00110000", -- 3      **
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11111110", -- 7    *******
    "11000000", -- 8    **
    "11000000", -- 9    **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x83
    "00000000", -- 0
    "00010000", -- 1       *
    "00111000", -- 2      ***
    "01101100", -- 3     ** **
    "00000000", -- 4
    "01111000", -- 5     ****
    "00001100", -- 6        **
    "01111100", -- 7     *****
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x84
    "00000000", -- 0
    "00000000", -- 1
    "11001100", -- 2    **  **
    "00000000", -- 3
    "00000000", -- 4
    "01111000", -- 5     ****
    "00001100", -- 6        **
    "01111100", -- 7     *****
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x85
    "00000000", -- 0
    "01100000", -- 1     **
    "00110000", -- 2      **
    "00011000", -- 3       **
    "00000000", -- 4
    "01111000", -- 5     ****
    "00001100", -- 6        **
    "01111100", -- 7     *****
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x86
    "00000000", -- 0
    "00111000", -- 1      ***
    "01101100", -- 2     ** **
    "00111000", -- 3      ***
    "00000000", -- 4
    "01111000", -- 5     ****
    "00001100", -- 6        **
    "01111100", -- 7     *****
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x87
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00111100", -- 4      ****
    "01100110", -- 5     **  **
    "01100000", -- 6     **
    "01100000", -- 7     **
    "01100110", -- 8     **  **
    "00111100", -- 9      ****
    "00001100", -- a        **
    "00000110", -- b         **
    "00111100", -- c      ****
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x88
    "00000000", -- 0
    "00010000", -- 1       *
    "00111000", -- 2      ***
    "01101100", -- 3     ** **
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11111110", -- 7    *******
    "11000000", -- 8    **
    "11000000", -- 9    **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x89
    "00000000", -- 0
    "00000000", -- 1
    "11000110", -- 2    **   **
    "00000000", -- 3
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11111110", -- 7    *******
    "11000000", -- 8    **
    "11000000", -- 9    **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x8A
    "00000000", -- 0
    "01100000", -- 1     **
    "00110000", -- 2      **
    "00011000", -- 3       **
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11111110", -- 7    *******
    "11000000", -- 8    **
    "11000000", -- 9    **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x8B
    "00000000", -- 0
    "00000000", -- 1
    "01100110", -- 2     **  **
    "00000000", -- 3
    "00000000", -- 4
    "00111000", -- 5      ***
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x8C
    "00000000", -- 0
    "00011000", -- 1       **
    "00111100", -- 2      ****
    "01100110", -- 3     **  **
    "00000000", -- 4
    "00111000", -- 5      ***
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x8D
    "00000000", -- 0
    "01100000", -- 1     **
    "00110000", -- 2      **
    "00011000", -- 3       **
    "00000000", -- 4
    "00111000", -- 5      ***
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x8E
    "00000000", -- 0
    "11000110", -- 1    **   **
    "00000000", -- 2
    "00010000", -- 3       *
    "00111000", -- 4      ***
    "01101100", -- 5     ** **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11111110", -- 8    *******
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "11000110", -- b    **   **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x8F
    "00111000", -- 0      ***
    "01101100", -- 1     ** **
    "00111000", -- 2      ***
    "00000000", -- 3
    "00111000", -- 4      ***
    "01101100", -- 5     ** **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11111110", -- 8    *******
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "11000110", -- b    **   **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x90
    "00011000", -- 0       **
    "00110000", -- 1      **
    "01100000", -- 2     **
    "00000000", -- 3
    "11111110", -- 4    *******
    "01100110", -- 5     **  **
    "01100000", -- 6     **
    "01111100", -- 7     *****
    "01100000", -- 8     **
    "01100000", -- 9     **
    "01100110", -- a     **  **
    "11111110", -- b    *******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x91
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01101110", -- 5     ** ***
    "00111011", -- 6      *** **
    "00011011", -- 7       ** **
    "01111110", -- 8     ******
    "11011000", -- 9    ** **
    "11011100", -- a    ** ***
    "01110111", -- b     *** ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x92
    "00000000", -- 0
    "00000000", -- 1
    "00111110", -- 2      *****
    "01101100", -- 3     ** **
    "11001100", -- 4    **  **
    "11001100", -- 5    **  **
    "11111110", -- 6    *******
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "11001110", -- b    **  ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x93
    "00000000", -- 0
    "00010000", -- 1       *
    "00111000", -- 2      ***
    "01101100", -- 3     ** **
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x94
    "00000000", -- 0
    "00000000", -- 1
    "11000110", -- 2    **   **
    "00000000", -- 3
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x95
    "00000000", -- 0
    "01100000", -- 1     **
    "00110000", -- 2      **
    "00011000", -- 3       **
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x96
    "00000000", -- 0
    "00110000", -- 1      **
    "01111000", -- 2     ****
    "11001100", -- 3    **  **
    "00000000", -- 4
    "11001100", -- 5    **  **
    "11001100", -- 6    **  **
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x97
    "00000000", -- 0
    "01100000", -- 1     **
    "00110000", -- 2      **
    "00011000", -- 3       **
    "00000000", -- 4
    "11001100", -- 5    **  **
    "11001100", -- 6    **  **
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x98
    "00000000", -- 0
    "00000000", -- 1
    "11000110", -- 2    **   **
    "00000000", -- 3
    "00000000", -- 4
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111110", -- b     ******
    "00000110", -- c         **
    "00001100", -- d        **
    "01111000", -- e     ****
    "00000000", -- f
    -- codigo x99
    "00000000", -- 0
    "11000110", -- 1    **   **
    "00000000", -- 2
    "01111100", -- 3     *****
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x9A
    "00000000", -- 0
    "11000110", -- 1    **   **
    "00000000", -- 2
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x9B
    "00000000", -- 0
    "00011000", -- 1       **
    "00011000", -- 2       **
    "01111110", -- 3     ******
    "11000011", -- 4    **    **
    "11000000", -- 5    **
    "11000000", -- 6    **
    "11000000", -- 7    **
    "11000011", -- 8    **    **
    "01111110", -- 9     ******
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x9C
    "00000000", -- 0
    "00111000", -- 1      ***
    "01101100", -- 2     ** **
    "01100100", -- 3     **  *
    "01100000", -- 4     **
    "11110000", -- 5    ****
    "01100000", -- 6     **
    "01100000", -- 7     **
    "01100000", -- 8     **
    "01100000", -- 9     **
    "11100110", -- a    ***  **
    "11111100", -- b    ******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x9D
    "00000000", -- 0
    "00000000", -- 1
    "11000011", -- 2    **    **
    "01100110", -- 3     **  **
    "00111100", -- 4      ****
    "00011000", -- 5       **
    "11111111", -- 6    ********
    "00011000", -- 7       **
    "11111111", -- 8    ********
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x9E
    "00000000", -- 0
    "11111100", -- 1    ******
    "01100110", -- 2     **  **
    "01100110", -- 3     **  **
    "01111100", -- 4     *****
    "01100010", -- 5     **   *
    "01100110", -- 6     **  **
    "01101111", -- 7     ** ****
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "11110011", -- b    ****  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo x9F
    "00000000", -- 0
    "00001110", -- 1        ***
    "00011011", -- 2       ** **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "01111110", -- 6     ******
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "11011000", -- c    ** **
    "01110000", -- d     ***
    "00000000", -- e
    "00000000", -- f
    -- codigo xA0
    "00000000", -- 0
    "00011000", -- 1       **
    "00110000", -- 2      **
    "01100000", -- 3     **
    "00000000", -- 4
    "01111000", -- 5     ****
    "00001100", -- 6        **
    "01111100", -- 7     *****
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xA1
    "00000000", -- 0
    "00001100", -- 1        **
    "00011000", -- 2       **
    "00110000", -- 3      **
    "00000000", -- 4
    "00111000", -- 5      ***
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xA2
    "00000000", -- 0
    "00011000", -- 1       **
    "00110000", -- 2      **
    "01100000", -- 3     **
    "00000000", -- 4
    "01111100", -- 5     *****
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xA3
    "00000000", -- 0
    "00011000", -- 1       **
    "00110000", -- 2      **
    "01100000", -- 3     **
    "00000000", -- 4
    "11001100", -- 5    **  **
    "11001100", -- 6    **  **
    "11001100", -- 7    **  **
    "11001100", -- 8    **  **
    "11001100", -- 9    **  **
    "11001100", -- a    **  **
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xA4
    "00000000", -- 0
    "00000000", -- 1
    "01110110", -- 2     *** **
    "11011100", -- 3    ** ***
    "00000000", -- 4
    "11011100", -- 5    ** ***
    "01100110", -- 6     **  **
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "01100110", -- b     **  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xA5
    "01110110", -- 0     *** **
    "11011100", -- 1    ** ***
    "00000000", -- 2
    "11000110", -- 3    **   **
    "11100110", -- 4    ***  **
    "11110110", -- 5    **** **
    "11111110", -- 6    *******
    "11011110", -- 7    ** ****
    "11001110", -- 8    **  ***
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "11000110", -- b    **   **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xA6
    "00000000", -- 0
    "00111100", -- 1      ****
    "01101100", -- 2     ** **
    "01101100", -- 3     ** **
    "00111110", -- 4      *****
    "00000000", -- 5
    "01111110", -- 6     ******
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xA7
    "00000000", -- 0
    "00111000", -- 1      ***
    "01101100", -- 2     ** **
    "01101100", -- 3     ** **
    "00111000", -- 4      ***
    "00000000", -- 5
    "01111100", -- 6     *****
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xA8
    "00000000", -- 0
    "00000000", -- 1
    "00110000", -- 2      **
    "00110000", -- 3      **
    "00000000", -- 4
    "00110000", -- 5      **
    "00110000", -- 6      **
    "01100000", -- 7     **
    "11000000", -- 8    **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "01111100", -- b     *****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xA9
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "11111110", -- 6    *******
    "11000000", -- 7    **
    "11000000", -- 8    **
    "11000000", -- 9    **
    "11000000", -- a    **
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xAA
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "11111110", -- 6    *******
    "00000110", -- 7         **
    "00000110", -- 8         **
    "00000110", -- 9         **
    "00000110", -- a         **
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xAB
    "00000000", -- 0
    "11000000", -- 1    **
    "11000000", -- 2    **
    "11000010", -- 3    **    *
    "11000110", -- 4    **   **
    "11001100", -- 5    **  **
    "00011000", -- 6       **
    "00110000", -- 7      **
    "01100000", -- 8     **
    "11001110", -- 9    **  ***
    "10011011", -- a    *  ** **
    "00000110", -- b         **
    "00001100", -- c        **
    "00011111", -- d       *****
    "00000000", -- e
    "00000000", -- f
    -- codigo xAC
    "00000000", -- 0
    "11000000", -- 1    **
    "11000000", -- 2    **
    "11000010", -- 3    **    *
    "11000110", -- 4    **   **
    "11001100", -- 5    **  **
    "00011000", -- 6       **
    "00110000", -- 7      **
    "01100110", -- 8     **  **
    "11001110", -- 9    **  ***
    "10010110", -- a    *  * **
    "00111110", -- b      *****
    "00000110", -- c         **
    "00000110", -- d         **
    "00000000", -- e
    "00000000", -- f
    -- codigo xAD
    "00000000", -- 0
    "00000000", -- 1
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00000000", -- 4
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00111100", -- 8      ****
    "00111100", -- 9      ****
    "00111100", -- a      ****
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xAE
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00110110", -- 5      ** **
    "01101100", -- 6     ** **
    "11011000", -- 7    ** **
    "01101100", -- 8     ** **
    "00110110", -- 9      ** **
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xAF
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11011000", -- 5    ** **
    "01101100", -- 6     ** **
    "00110110", -- 7      ** **
    "01101100", -- 8     ** **
    "11011000", -- 9    ** **
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xB0
    "00010001", -- 0       *   *
    "01000100", -- 1     *   *
    "00010001", -- 2       *   *
    "01000100", -- 3     *   *
    "00010001", -- 4       *   *
    "01000100", -- 5     *   *
    "00010001", -- 6       *   *
    "01000100", -- 7     *   *
    "00010001", -- 8       *   *
    "01000100", -- 9     *   *
    "00010001", -- a       *   *
    "01000100", -- b     *   *
    "00010001", -- c       *   *
    "01000100", -- d     *   *
    "00010001", -- e       *   *
    "01000100", -- f     *   *
    -- codigo xB1
    "01010101", -- 0     * * * *
    "10101010", -- 1    * * * *
    "01010101", -- 2     * * * *
    "10101010", -- 3    * * * *
    "01010101", -- 4     * * * *
    "10101010", -- 5    * * * *
    "01010101", -- 6     * * * *
    "10101010", -- 7    * * * *
    "01010101", -- 8     * * * *
    "10101010", -- 9    * * * *
    "01010101", -- a     * * * *
    "10101010", -- b    * * * *
    "01010101", -- c     * * * *
    "10101010", -- d    * * * *
    "01010101", -- e     * * * *
    "10101010", -- f    * * * *
    -- codigo xB2
    "11011101", -- 0    ** *** *
    "01110111", -- 1     *** ***
    "11011101", -- 2    ** *** *
    "01110111", -- 3     *** ***
    "11011101", -- 4    ** *** *
    "01110111", -- 5     *** ***
    "11011101", -- 6    ** *** *
    "01110111", -- 7     *** ***
    "11011101", -- 8    ** *** *
    "01110111", -- 9     *** ***
    "11011101", -- a    ** *** *
    "01110111", -- b     *** ***
    "11011101", -- c    ** *** *
    "01110111", -- d     *** ***
    "11011101", -- e    ** *** *
    "01110111", -- f     *** ***
    -- codigo xB3
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xB4
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "11111000", -- 7    *****
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xB5
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "11111000", -- 5    *****
    "00011000", -- 6       **
    "11111000", -- 7    *****
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xB6
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "00110110", -- 5      ** **
    "00110110", -- 6      ** **
    "11110110", -- 7    **** **
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xB7
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "11111110", -- 7    *******
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xB8
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11111000", -- 5    *****
    "00011000", -- 6       **
    "11111000", -- 7    *****
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xB9
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "11110110", -- 5    **** **
    "00000110", -- 6         **
    "11110110", -- 7    **** **
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xBA
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "00110110", -- 5      ** **
    "00110110", -- 6      ** **
    "00110110", -- 7      ** **
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xBB
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11111110", -- 5    *******
    "00000110", -- 6         **
    "11110110", -- 7    **** **
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xBC
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "11110110", -- 5    **** **
    "00000110", -- 6         **
    "11111110", -- 7    *******
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xBD
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "00110110", -- 5      ** **
    "00110110", -- 6      ** **
    "11111110", -- 7    *******
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xBE
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "11111000", -- 5    *****
    "00011000", -- 6       **
    "11111000", -- 7    *****
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xBF
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "11111000", -- 7    *****
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xC0
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011111", -- 7       *****
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xC1
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "11111111", -- 7    ********
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xC2
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "11111111", -- 7    ********
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xC3
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011111", -- 7       *****
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xC4
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "11111111", -- 7    ********
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xC5
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "11111111", -- 7    ********
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xC6
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011111", -- 5       *****
    "00011000", -- 6       **
    "00011111", -- 7       *****
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xC7
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "00110110", -- 5      ** **
    "00110110", -- 6      ** **
    "00110111", -- 7      ** ***
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xC8
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "00110111", -- 5      ** ***
    "00110000", -- 6      **
    "00111111", -- 7      ******
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xC9
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00111111", -- 5      ******
    "00110000", -- 6      **
    "00110111", -- 7      ** ***
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xCA
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "11110111", -- 5    **** ***
    "00000000", -- 6
    "11111111", -- 7    ********
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xCB
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11111111", -- 5    ********
    "00000000", -- 6
    "11110111", -- 7    **** ***
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xCC
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "00110111", -- 5      ** ***
    "00110000", -- 6      **
    "00110111", -- 7      ** ***
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xCD
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11111111", -- 5    ********
    "00000000", -- 6
    "11111111", -- 7    ********
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xCE
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "11110111", -- 5    **** ***
    "00000000", -- 6
    "11110111", -- 7    **** ***
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xCF
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "11111111", -- 5    ********
    "00000000", -- 6
    "11111111", -- 7    ********
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xD0
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "00110110", -- 5      ** **
    "00110110", -- 6      ** **
    "11111111", -- 7    ********
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xD1
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "11111111", -- 5    ********
    "00000000", -- 6
    "11111111", -- 7    ********
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xD2
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "11111111", -- 7    ********
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xD3
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "00110110", -- 5      ** **
    "00110110", -- 6      ** **
    "00111111", -- 7      ******
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xD4
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011111", -- 5       *****
    "00011000", -- 6       **
    "00011111", -- 7       *****
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xD5
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00011111", -- 5       *****
    "00011000", -- 6       **
    "00011111", -- 7       *****
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xD6
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00111111", -- 7      ******
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xD7
    "00110110", -- 0      ** **
    "00110110", -- 1      ** **
    "00110110", -- 2      ** **
    "00110110", -- 3      ** **
    "00110110", -- 4      ** **
    "00110110", -- 5      ** **
    "00110110", -- 6      ** **
    "11111111", -- 7    ********
    "00110110", -- 8      ** **
    "00110110", -- 9      ** **
    "00110110", -- a      ** **
    "00110110", -- b      ** **
    "00110110", -- c      ** **
    "00110110", -- d      ** **
    "00110110", -- e      ** **
    "00110110", -- f      ** **
    -- codigo xD8
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "11111111", -- 5    ********
    "00011000", -- 6       **
    "11111111", -- 7    ********
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xD9
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "11111000", -- 7    *****
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xDA
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00011111", -- 7       *****
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xDB
    "11111111", -- 0    ********
    "11111111", -- 1    ********
    "11111111", -- 2    ********
    "11111111", -- 3    ********
    "11111111", -- 4    ********
    "11111111", -- 5    ********
    "11111111", -- 6    ********
    "11111111", -- 7    ********
    "11111111", -- 8    ********
    "11111111", -- 9    ********
    "11111111", -- a    ********
    "11111111", -- b    ********
    "11111111", -- c    ********
    "11111111", -- d    ********
    "11111111", -- e    ********
    "11111111", -- f    ********
    -- codigo xDC
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "11111111", -- 7    ********
    "11111111", -- 8    ********
    "11111111", -- 9    ********
    "11111111", -- a    ********
    "11111111", -- b    ********
    "11111111", -- c    ********
    "11111111", -- d    ********
    "11111111", -- e    ********
    "11111111", -- f    ********
    -- codigo xDD
    "11110000", -- 0    ****
    "11110000", -- 1    ****
    "11110000", -- 2    ****
    "11110000", -- 3    ****
    "11110000", -- 4    ****
    "11110000", -- 5    ****
    "11110000", -- 6    ****
    "11110000", -- 7    ****
    "11110000", -- 8    ****
    "11110000", -- 9    ****
    "11110000", -- a    ****
    "11110000", -- b    ****
    "11110000", -- c    ****
    "11110000", -- d    ****
    "11110000", -- e    ****
    "11110000", -- f    ****
    -- codigo xDE
    "00001111", -- 0        ****
    "00001111", -- 1        ****
    "00001111", -- 2        ****
    "00001111", -- 3        ****
    "00001111", -- 4        ****
    "00001111", -- 5        ****
    "00001111", -- 6        ****
    "00001111", -- 7        ****
    "00001111", -- 8        ****
    "00001111", -- 9        ****
    "00001111", -- a        ****
    "00001111", -- b        ****
    "00001111", -- c        ****
    "00001111", -- d        ****
    "00001111", -- e        ****
    "00001111", -- f        ****
    -- codigo xDF
    "11111111", -- 0    ********
    "11111111", -- 1    ********
    "11111111", -- 2    ********
    "11111111", -- 3    ********
    "11111111", -- 4    ********
    "11111111", -- 5    ********
    "11111111", -- 6    ********
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE0
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01110110", -- 5     *** **
    "11011100", -- 6    ** ***
    "11011000", -- 7    ** **
    "11011000", -- 8    ** **
    "11011000", -- 9    ** **
    "11011100", -- a    ** ***
    "01110110", -- b     *** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE1
    "00000000", -- 0
    "00000000", -- 1
    "01111000", -- 2     ****
    "11001100", -- 3    **  **
    "11001100", -- 4    **  **
    "11001100", -- 5    **  **
    "11011000", -- 6    ** **
    "11001100", -- 7    **  **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "11001100", -- b    **  **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE2
    "00000000", -- 0
    "00000000", -- 1
    "11111110", -- 2    *******
    "11000110", -- 3    **   **
    "11000110", -- 4    **   **
    "11000000", -- 5    **
    "11000000", -- 6    **
    "11000000", -- 7    **
    "11000000", -- 8    **
    "11000000", -- 9    **
    "11000000", -- a    **
    "11000000", -- b    **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE3
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "11111110", -- 4    *******
    "01101100", -- 5     ** **
    "01101100", -- 6     ** **
    "01101100", -- 7     ** **
    "01101100", -- 8     ** **
    "01101100", -- 9     ** **
    "01101100", -- a     ** **
    "01101100", -- b     ** **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE4
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "11111110", -- 3    *******
    "11000110", -- 4    **   **
    "01100000", -- 5     **
    "00110000", -- 6      **
    "00011000", -- 7       **
    "00110000", -- 8      **
    "01100000", -- 9     **
    "11000110", -- a    **   **
    "11111110", -- b    *******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE5
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01111110", -- 5     ******
    "11011000", -- 6    ** **
    "11011000", -- 7    ** **
    "11011000", -- 8    ** **
    "11011000", -- 9    ** **
    "11011000", -- a    ** **
    "01110000", -- b     ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE6
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "01100110", -- 4     **  **
    "01100110", -- 5     **  **
    "01100110", -- 6     **  **
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "01111100", -- 9     *****
    "01100000", -- a     **
    "01100000", -- b     **
    "11000000", -- c    **
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE7
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "01110110", -- 4     *** **
    "11011100", -- 5    ** ***
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE8
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "01111110", -- 3     ******
    "00011000", -- 4       **
    "00111100", -- 5      ****
    "01100110", -- 6     **  **
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "00111100", -- 9      ****
    "00011000", -- a       **
    "01111110", -- b     ******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xE9
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00111000", -- 3      ***
    "01101100", -- 4     ** **
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11111110", -- 7    *******
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "01101100", -- a     ** **
    "00111000", -- b      ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xEA
    "00000000", -- 0
    "00000000", -- 1
    "00111000", -- 2      ***
    "01101100", -- 3     ** **
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "01101100", -- 7     ** **
    "01101100", -- 8     ** **
    "01101100", -- 9     ** **
    "01101100", -- a     ** **
    "11101110", -- b    *** ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xEB
    "00000000", -- 0
    "00000000", -- 1
    "00011110", -- 2       ****
    "00110000", -- 3      **
    "00011000", -- 4       **
    "00001100", -- 5        **
    "00111110", -- 6      *****
    "01100110", -- 7     **  **
    "01100110", -- 8     **  **
    "01100110", -- 9     **  **
    "01100110", -- a     **  **
    "00111100", -- b      ****
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xEC
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01111110", -- 5     ******
    "11011011", -- 6    ** ** **
    "11011011", -- 7    ** ** **
    "11011011", -- 8    ** ** **
    "01111110", -- 9     ******
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xED
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000011", -- 3          **
    "00000110", -- 4         **
    "01111110", -- 5     ******
    "11011011", -- 6    ** ** **
    "11011011", -- 7    ** ** **
    "11110011", -- 8    ****  **
    "01111110", -- 9     ******
    "01100000", -- a     **
    "11000000", -- b    **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xEE
    "00000000", -- 0
    "00000000", -- 1
    "00011100", -- 2       ***
    "00110000", -- 3      **
    "01100000", -- 4     **
    "01100000", -- 5     **
    "01111100", -- 6     *****
    "01100000", -- 7     **
    "01100000", -- 8     **
    "01100000", -- 9     **
    "00110000", -- a      **
    "00011100", -- b       ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xEF
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "01111100", -- 3     *****
    "11000110", -- 4    **   **
    "11000110", -- 5    **   **
    "11000110", -- 6    **   **
    "11000110", -- 7    **   **
    "11000110", -- 8    **   **
    "11000110", -- 9    **   **
    "11000110", -- a    **   **
    "11000110", -- b    **   **
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xF0
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "11111110", -- 4    *******
    "00000000", -- 5
    "00000000", -- 6
    "11111110", -- 7    *******
    "00000000", -- 8
    "00000000", -- 9
    "11111110", -- a    *******
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xF1
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00011000", -- 4       **
    "00011000", -- 5       **
    "01111110", -- 6     ******
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00000000", -- 9
    "00000000", -- a
    "11111111", -- b    ********
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xF2
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00110000", -- 3      **
    "00011000", -- 4       **
    "00001100", -- 5        **
    "00000110", -- 6         **
    "00001100", -- 7        **
    "00011000", -- 8       **
    "00110000", -- 9      **
    "00000000", -- a
    "01111110", -- b     ******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xF3
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00001100", -- 3        **
    "00011000", -- 4       **
    "00110000", -- 5      **
    "01100000", -- 6     **
    "00110000", -- 7      **
    "00011000", -- 8       **
    "00001100", -- 9        **
    "00000000", -- a
    "01111110", -- b     ******
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xF4
    "00000000", -- 0
    "00000000", -- 1
    "00001110", -- 2        ***
    "00011011", -- 3       ** **
    "00011011", -- 4       ** **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00011000", -- 9       **
    "00011000", -- a       **
    "00011000", -- b       **
    "00011000", -- c       **
    "00011000", -- d       **
    "00011000", -- e       **
    "00011000", -- f       **
    -- codigo xF5
    "00011000", -- 0       **
    "00011000", -- 1       **
    "00011000", -- 2       **
    "00011000", -- 3       **
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00011000", -- 6       **
    "00011000", -- 7       **
    "11011000", -- 8    ** **
    "11011000", -- 9    ** **
    "11011000", -- a    ** **
    "01110000", -- b     ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xF6
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00011000", -- 4       **
    "00011000", -- 5       **
    "00000000", -- 6
    "01111110", -- 7     ******
    "00000000", -- 8
    "00011000", -- 9       **
    "00011000", -- a       **
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xF7
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "01110110", -- 5     *** **
    "11011100", -- 6    ** ***
    "00000000", -- 7
    "01110110", -- 8     *** **
    "11011100", -- 9    ** ***
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xF8
    "00000000", -- 0
    "00111000", -- 1      ***
    "01101100", -- 2     ** **
    "01101100", -- 3     ** **
    "00111000", -- 4      ***
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xF9
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00011000", -- 7       **
    "00011000", -- 8       **
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xFA
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00011000", -- 8       **
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xFB
    "00000000", -- 0
    "00001111", -- 1        ****
    "00001100", -- 2        **
    "00001100", -- 3        **
    "00001100", -- 4        **
    "00001100", -- 5        **
    "00001100", -- 6        **
    "11101100", -- 7    *** **
    "01101100", -- 8     ** **
    "01101100", -- 9     ** **
    "00111100", -- a      ****
    "00011100", -- b       ***
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xFC
    "00000000", -- 0
    "11011000", -- 1    ** **
    "01101100", -- 2     ** **
    "01101100", -- 3     ** **
    "01101100", -- 4     ** **
    "01101100", -- 5     ** **
    "01101100", -- 6     ** **
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xFD
    "00000000", -- 0
    "01110000", -- 1     ***
    "11011000", -- 2    ** **
    "00110000", -- 3      **
    "01100000", -- 4     **
    "11001000", -- 5    **  *
    "11111000", -- 6    *****
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xFE
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "01111100", -- 4     *****
    "01111100", -- 5     *****
    "01111100", -- 6     *****
    "01111100", -- 7     *****
    "01111100", -- 8     *****
    "01111100", -- 9     *****
    "01111100", -- a     *****
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000", -- f
    -- codigo xFF
    "00000000", -- 0
    "00000000", -- 1
    "00000000", -- 2
    "00000000", -- 3
    "00000000", -- 4
    "00000000", -- 5
    "00000000", -- 6
    "00000000", -- 7
    "00000000", -- 8
    "00000000", -- 9
    "00000000", -- a
    "00000000", -- b
    "00000000", -- c
    "00000000", -- d
    "00000000", -- e
    "00000000"  -- f
  );

begin

  -- addr register to infer block RAM
  --   process (clk)
  --   begin
  --      if (clk'event and clk = '1') then
  addr_reg <= addr;
  --      end if;
  --   end process;
  data <= ROM(to_integer(unsigned(addr_reg)));

end architecture vga_font_rom_arch;

